>A, Ala, Alanine
GCT
GCC
GCA
GCG
>D, Asp, Aspartic acid
GAT
GAC
>F, Phe, Phenylalanine
TTT
TTC
>H, His, Histidine
CAT
CAC
>K, Lys, Lysine
AAA
AAG
>M, Met, Methionine
ATG
>P, Pro, Proline
CCT
CCC
CCA
CCG
>R, Arg, Arginine
CGT
CGC
CGA
CGG
AGA
AGG
>T, Thr, Threonine
ACT
ACC
ACA
ACG
>W, Trp, Tryptophan
TGG
>C, Cys, Cysteine
TGT
TGC
>E, Glu, Glutamic Acid
GAA
GAG
>G, Gly, Glycine
GGT
GGC
GGA
GGG
>I, Ile, Isoleucine
ATT
ATC
ATA
>L, Leu, Leucine
TTA
TTG
CTT
CTC
CTA
CTG
>N, Asn, Asparagine
AAT
AAC
>Q, Gln, Glutamine
CAA
CAG
>S, Ser, Serine
TCT
TCC
TCA
TCG
AGT
AGC
>V, Val, Valine
GTT
GTC
GTA
GTG
>Y, Tyr, Tyrosine
TAT
TAC
